class read_xtn extends uvm_sequence_item;
`uvm_object_utils(read_xtn)

function new(string name="read_xtn");
super.new(name);
endfunction

endclass

