class wr_agt_config extends uvm_object;
`uvm_object_utils(wr_agt_config)

virtual fifo_if vif;

function new(string name="wr_agt_config");
super.new(name);
endfunction

uvm_active_passive_enum is_active=UVM_ACTIVE;

endclass
