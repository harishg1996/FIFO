class rd_agt_sequencer extends uvm_sequencer#(read_xtn);
`uvm_component_utils(rd_agt_sequencer)

function new(string name="rd_agt_sequencer",uvm_component parent);
super.new(name,parent);
endfunction

endclass

